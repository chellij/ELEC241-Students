entity task2p1 is

	port
	(
		-- Input ports
		X	: in  bit;

		-- Output ports
		Y	: out bit
	);
end task2p1;



-- Library Clause(s) (optional)
-- Use Clause(s) (optional)

architecture task2p1_v1 of task2p1 is

	-- Declarations (optional)

begin

	Y <= ;

end task2p1_v1;
